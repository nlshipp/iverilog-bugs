/*******************************************************************************
* Copyright 2009, Cypress Semiconductor Corporation.  All rights reserved.
* You may use this file only in accordance with the license, terms, conditions, 
* disclaimers, and limitations in the end user license agreement accompanying 
* the software package with which this file was provided.
********************************************************************************/

//
//	PSoC3 RTL Components
//

`ifdef PSOC3_RTL_ALREADY_INCLUDED
    // Only include the rest of this file once.
`else
`define PSOC3_RTL_ALREADY_INCLUDED
`define TRUE  1
`define FALSE 0

//
//	cy_psoc3_dp
//

`include "cy_psoc3_dp.v"

//
// 	cy_psoc3_carry
//

module cy_psoc3_carry (cin, cpt0, cpt1, sum, cout);
    input	cin;
    input	cpt0;
    input	cpt1;
    output	sum;
    output	cout;

    wire sum	= (cpt0 | cpt1) ^~ cin;
    wire cout	= (~cin & cpt0) | (cin & ~cpt1);
endmodule

//
//	cy_psoc3_control
//

module cy_psoc3_control (reset, clock, control);
    input		reset;
    input		clock;
    output	[07:00]	control;

    parameter	[07:00]	cy_init_value	= 8'b0;
    parameter		cy_force_order	= `FALSE;
    parameter		cy_ext_reset	= `FALSE;
    parameter	[07:00]	cy_ctrl_mode_1	= 8'b0;
    parameter	[07:00]	cy_ctrl_mode_0	= 8'b0;

    reg		[07:00] cpu_control;
    reg		[07:00] syn_control;
    reg		[07:00]	cpu_data;
    reg			cpu_write;
    reg			cpu_clock;	// Generated by the test bench.

    initial cpu_control = cy_init_value;

    // Synchronous reset
    reg [07:00] sync_reset;
    always @(posedge clock)
    begin
    	sync_reset = cy_ctrl_mode_1 & syn_control;
    end

    // The original Control Register
    always @(posedge reset or posedge (| sync_reset) or posedge cpu_write)
    begin
    	if (reset && cy_ext_reset)
	    cpu_control <= 8'b0;
	else if (sync_reset)
	    cpu_control <= cpu_control & ~sync_reset;
	else if (cpu_write)
	    cpu_control <= cpu_data;
    end

    // Generate the synchronizing FFs
    always @(posedge clock or posedge reset or posedge (| sync_reset))
    begin
	if (reset)
	    syn_control <= 8'b0;
	else if (sync_reset)
	    syn_control <= syn_control & ~sync_reset;
	else
	    syn_control <= cpu_control;
    end

    wire [07:00] control = ( cy_ctrl_mode_0 & syn_control) |
			   (~cy_ctrl_mode_0 & cpu_control);

    // Task to write the control register via the CPU.
    task control_write;
    	input [07:00] data;
    begin
	cpu_data = data;
    	@(posedge cpu_clock)
	cpu_write <= 1'b1;
	@(posedge cpu_clock)
	cpu_write <= 1'b0;
    end
    endtask

endmodule

//
//	cy_psoc3_status w/o interrupt
//

module cy_psoc3_status (reset, clock, status);
    input		reset;
    input		clock;
    input	[07:00]	status;

    parameter		cy_force_order	= `FALSE;
    parameter	[07:00]	cy_md_select	= 8'b00000000;

    reg			cpu_clock;		// Generated by the test bench.
    reg			read_sig = 0;		// Trigger the reset_on_read.
    reg			reset_on_read = 0;	// Clears register on CPU read.

    reg [07:00] status_reg;
    always @(posedge clock or posedge reset or posedge reset_on_read)
    begin
	if (reset || reset_on_read)
	    status_reg <= 0;
	else
	    status_reg <=  status | status_reg;
    end

    reg [07:00] status_to_cpu;
    always @(status or status_reg)
    begin
	status_to_cpu[0] <= cy_md_select[0] ? status_reg[0] : status[0];
	status_to_cpu[1] <= cy_md_select[1] ? status_reg[1] : status[1];
	status_to_cpu[2] <= cy_md_select[2] ? status_reg[2] : status[2];
	status_to_cpu[3] <= cy_md_select[3] ? status_reg[3] : status[3];
	status_to_cpu[4] <= cy_md_select[4] ? status_reg[4] : status[4];
	status_to_cpu[5] <= cy_md_select[5] ? status_reg[5] : status[5];
	status_to_cpu[6] <= cy_md_select[6] ? status_reg[6] : status[6];
	status_to_cpu[7] <= cy_md_select[7] ? status_reg[7] : status[7];
    end

    // Reset the status register if a CPU read has occurred.
    always @(posedge read_sig)
    begin
    	@(posedge cpu_clock)
	reset_on_read <= 1'b1;
	@(posedge cpu_clock)
	reset_on_read <= 1'b0;
    end

    // Read the status register via the CPU (and start the reset_on_read).
    task status_read;
    	output [07:00] data;
    begin
	data <= status_to_cpu;
	read_sig <= 1;
	# 1;
	read_sig <= 0;
    end
    endtask

endmodule

//
//	cy_psoc3_status with interrupt
//

module cy_psoc3_statusi (reset, clock, status, interrupt);
    input		reset;
    input		clock;
    input	[06:00]	status;
    output		interrupt;

    parameter		cy_force_order	= `FALSE;
    parameter	[06:00]	cy_md_select	= 7'b0000000;
    parameter	[06:00]	cy_int_mask	= 7'b0000000;

    reg			cpu_clock;		// Generated by the test bench.
    reg			read_sig = 0;		// Trigger the reset_on_read.
    reg			reset_on_read = 0;	// Clears register on CPU read.

    // Instantiate Virtual Auxilliary Control & Mask Registers for MCU accesses
    reg 		actl;
    reg		[06:00]	mask;
    wire		int_en = actl;
    initial
    begin
	actl = 1'b1;
	mask = cy_int_mask;
    end

    reg [06:00] status_reg;
    always @(posedge clock or posedge reset or posedge reset_on_read)
    begin
    	if (reset || reset_on_read)
	    status_reg <= 0;
	else
	    status_reg <= status | status_reg;
    end

    reg [06:00] status_to_cpu;		// Available to the CPU
    always @(status or status_reg)
    begin
	status_to_cpu[0] <= cy_md_select[0] ? status_reg[0] : status[0];
	status_to_cpu[1] <= cy_md_select[1] ? status_reg[1] : status[1];
	status_to_cpu[2] <= cy_md_select[2] ? status_reg[2] : status[2];
	status_to_cpu[3] <= cy_md_select[3] ? status_reg[3] : status[3];
	status_to_cpu[4] <= cy_md_select[4] ? status_reg[4] : status[4];
	status_to_cpu[5] <= cy_md_select[5] ? status_reg[5] : status[5];
	status_to_cpu[6] <= cy_md_select[6] ? status_reg[6] : status[6];
    end

    assign interrupt = |(mask & status_to_cpu) & int_en;

    // Reset the statusi register if a CPU read has occurred.
    always @(posedge read_sig)
    begin
    	@(posedge cpu_clock)
	reset_on_read <= 1'b1;
	@(posedge cpu_clock)
	reset_on_read <= 1'b0;
    end

    // Read the statusi register via the CPU (and start the reset_on_read).
    task status_read;
    	output [06:00] data;
    begin
	data <= status_to_cpu;
	read_sig <= 1;
	# 1;
	read_sig <= 0;
    end
    endtask

endmodule

//
//	cy_psoc3_sync
//

module cy_psoc3_sync (clock, sc_in, sc_out);

    input	clock;
    input 	sc_in;
    output	sc_out;

    reg	 s_reg  = 1'b0;
    reg  sc_out = 1'b0;
    always @(posedge clock)
    begin
    	s_reg  <= sc_in;
	sc_out <= s_reg;
    end

endmodule


//
//	cy_psoc3_udb_clock_enable_v1_0
//

module cy_psoc3_udb_clock_enable_v1_0 (clock_in, enable, clock_out);

    input	clock_in;
    input	enable;
    output	clock_out;

    parameter	sync_mode = `FALSE;

    wire clock_out = (sync_mode == `FALSE) ? enable  & clock_in :
					    (enable) ? clock_in : 1'b0;

endmodule

//
//	cy_isr_v1_0
//

module cy_isr_v1_0 (int_signal);
    input		int_signal;
endmodule

//
//	cy_dma_v1_0
//

module cy_dma_v1_0 (drq, trq, nrq);
    input		drq;
    input		trq;
    output		nrq;

    parameter		num_tds	= 0;
endmodule

//
//	cy_psoc3_count7
//

module cy_psoc3_count7 (clock, reset, load, enable, count, tc);
    input		clock;
    input		reset;
    input		load;
    input		enable;
    output	[06:00]	count;
    output		tc;

    parameter	[06:00]	cy_period	= 7'b1111111;
    parameter	[06:00]	cy_init_value	= 7'b0000000;
    parameter		cy_route_ld	= `FALSE;
    parameter		cy_route_en	= `FALSE;
    parameter		cy_alt_mode	= `FALSE;

    wire #0 clk = clock;

    // Instantiate a Virtual Auxilliary Control Register for MCU accesses
    reg 		actl;
    wire		count_start = actl;
    initial actl = 1'b1;

    // Power-on reset
    reg reset_sys;
    initial 
    begin
      reset_sys = 1'b0;
      #1;
      reset_sys = 1'b1;
      #1;
      reset_sys = 1'b0;
    end

    wire reset_blk = reset_sys | reset;

    // Simulate the 7-bit counter
    reg	[06:00] count;
    reg	[06:00] period_reg;
    wire	zero_detect;
    wire	real_load   = (cy_alt_mode)
			    ? zero_detect | (load &    enable)
			    : zero_detect | (load &   (cy_route_ld == `TRUE));
    wire	real_enable = (cy_alt_mode)
			    ? count_start &  enable
			    : count_start & (enable | (cy_route_en == `FALSE));

    initial period_reg <= cy_period;

    reg count_clk_en;
    always @(clk or real_enable)
    begin
	if (!clk)
	    count_clk_en <= real_enable;
    end
    wire count_clk = count_clk_en & clk;

    always @(posedge count_clk or posedge reset_blk)
    begin
	if (reset_blk)
	    count <= cy_init_value;
	else if (real_load)
	    count <= period_reg;
	else
	    count <= count - 1;
    end

    // Has the count reached 0?
    assign zero_detect = (count == 7'b0);

    // Registered terminal count
    reg tc_reg = 0;
    always @(posedge count_clk or posedge reset_blk)
    begin
      if (reset_blk)
	  tc_reg <= 1'b0;
      else
	  tc_reg <= zero_detect;
    end

    wire tc = (cy_alt_mode) ? (zero_detect & count_start) : tc_reg;

endmodule

//
//	cy_psoc3_dp8
//

module cy_psoc3_dp8 (reset, clk,
    cs_addr, route_si, route_ci, f0_load, f1_load, d0_load, d1_load,
    ce0, cl0, z0, ff0, ce1, cl1, z1, ff1, ov_msb, co_msb, cmsb, so,
    f0_bus_stat, f0_blk_stat, f1_bus_stat, f1_blk_stat,
    ce0_reg, cl0_reg, z0_reg, ff0_reg, ce1_reg, cl1_reg, z1_reg,
    ff1_reg, ov_msb_reg, co_msb_reg, cmsb_reg, so_reg,
    f0_bus_stat_reg, f0_blk_stat_reg, f1_bus_stat_reg, f1_blk_stat_reg);
    input		reset;
    input		clk;
    input	[02:00]	cs_addr;
    input		route_si;
    input		route_ci;
    input		f0_load;
    input		f1_load;
    input		d0_load;
    input		d1_load;
    output		ce0;
    output		cl0;
    output		z0;
    output		ff0;
    output		ce1;
    output		cl1;
    output		z1;
    output		ff1;
    output		ov_msb;
    output		co_msb;
    output		cmsb;
    output		so;
    output		f0_bus_stat;
    output		f0_blk_stat;
    output		f1_bus_stat;
    output		f1_blk_stat;
    output		ce0_reg;
    output		cl0_reg;
    output		z0_reg;
    output		ff0_reg;
    output		ce1_reg;
    output		cl1_reg;
    output		z1_reg;
    output		ff1_reg;
    output		ov_msb_reg;
    output		co_msb_reg;
    output		cmsb_reg;
    output		so_reg;
    output		f0_bus_stat_reg;
    output		f0_blk_stat_reg;
    output		f1_bus_stat_reg;
    output		f1_blk_stat_reg;

    parameter	[207:0] cy_dpconfig_a	= {128'h0,32'hFF00_FFFF,48'h0};
    parameter	[07:00] d0_init_a	= 8'b0;
    parameter	[07:00] d1_init_a	= 8'b0;
    parameter	[07:00] a0_init_a	= 8'b0;
    parameter	[07:00] a1_init_a	= 8'b0;
    parameter		ce0_sync	= 1'b1;
    parameter		cl0_sync	= 1'b1;
    parameter		z0_sync		= 1'b1;
    parameter		ff0_sync	= 1'b1;
    parameter		ce1_sync	= 1'b1;
    parameter		cl1_sync	= 1'b1;
    parameter		z1_sync		= 1'b1;
    parameter		ff1_sync	= 1'b1;
    parameter		ov_msb_sync	= 1'b1;
    parameter		co_msb_sync	= 1'b1;
    parameter		cmsb_sync	= 1'b1;
    parameter		so_sync		= 1'b1;
    parameter		f0_bus_sync	= 1'b1;
    parameter		f0_blk_sync	= 1'b1;
    parameter		f1_bus_sync	= 1'b1;
    parameter		f1_blk_sync	= 1'b1;

    defparam U0.cy_dpconfig	= cy_dpconfig_a;
    defparam U0.d0_init		= d0_init_a;
    defparam U0.d1_init		= d1_init_a;
    defparam U0.a0_init		= a0_init_a;
    defparam U0.a1_init		= a1_init_a;
    defparam U0.ce0_sync	= ce0_sync;
    defparam U0.cl0_sync	= cl0_sync;
    defparam U0.z0_sync		= z0_sync;
    defparam U0.ff0_sync	= ff0_sync;
    defparam U0.ce1_sync	= ce1_sync;
    defparam U0.cl1_sync	= cl1_sync;
    defparam U0.z1_sync		= z1_sync;
    defparam U0.ff1_sync	= ff1_sync;
    defparam U0.ov_msb_sync	= ov_msb_sync;
    defparam U0.co_msb_sync	= co_msb_sync;
    defparam U0.cmsb_sync	= cmsb_sync;
    defparam U0.so_sync		= so_sync;
    defparam U0.f0_bus_sync	= f0_bus_sync;
    defparam U0.f0_blk_sync	= f0_blk_sync;
    defparam U0.f1_bus_sync	= f1_bus_sync;
    defparam U0.f1_blk_sync	= f1_blk_sync;
    cy_psoc3_dp U0 (
	.reset			(reset),
	.clk			(clk),
	.cs_addr		(cs_addr),
	.route_si		(route_si),
	.route_ci		(route_ci),
	.f0_load		(f0_load),
	.f1_load		(f1_load),
	.d0_load		(d0_load),
	.d1_load		(d1_load),
	.ce0			(ce0),
	.cl0			(cl0),
	.z0			(z0),
	.ff0			(ff0),
	.ce1			(ce1),
	.cl1			(cl1),
	.z1			(z1),
	.ff1			(ff1),
	.ov_msb			(ov_msb),
	.co_msb			(co_msb),
	.cmsb			(cmsb),
	.so			(so),
	.f0_bus_stat		(f0_bus_stat),
	.f0_blk_stat		(f0_blk_stat),
	.f1_bus_stat		(f1_bus_stat),
	.f1_blk_stat		(f1_blk_stat),
	.ce0_reg		(ce0_reg),
	.cl0_reg		(cl0_reg),
	.z0_reg			(z0_reg),
	.ff0_reg		(ff0_reg),
	.ce1_reg		(ce1_reg),
	.cl1_reg		(cl1_reg),
	.z1_reg			(z1_reg),
	.ff1_reg		(ff1_reg),
	.ov_msb_reg		(ov_msb_reg),
	.co_msb_reg		(co_msb_reg),
	.cmsb_reg		(cmsb_reg),
	.so_reg			(so_reg),
	.f0_bus_stat_reg	(f0_bus_stat_reg),
	.f0_blk_stat_reg	(f0_blk_stat_reg),
	.f1_bus_stat_reg	(f1_bus_stat_reg),
	.f1_blk_stat_reg	(f1_blk_stat_reg),
	.ci			(1'b0),
	.co			(),
	.sir			(1'b0),
	.sor			(),
	.sil			(1'b0),
	.sol			(),
	.msbi			(1'b0),
	.msbo			(),
	.cei			(2'b00),
	.ceo			(),
	.cli			(2'b00),
	.clo			(),
	.zi			(2'b00),
	.zo			(),
	.fi			(2'b00),
	.fo			(),
	.capi			(2'b00),
	.capo			(),
	.cfbi			(1'b1),
	.cfbo			(),
	.pi			(8'b00000000),
	.po			());
endmodule

//
//	cy_psoc3_dp16
//

module cy_psoc3_dp16 (reset, clk,
    cs_addr, route_si, route_ci, f0_load, f1_load, d0_load, d1_load,
    ce0, cl0, z0, ff0, ce1, cl1, z1, ff1, ov_msb, co_msb, cmsb, so,
    f0_bus_stat, f0_blk_stat, f1_bus_stat, f1_blk_stat,
    ce0_reg, cl0_reg, z0_reg, ff0_reg, ce1_reg, cl1_reg, z1_reg,
    ff1_reg, ov_msb_reg, co_msb_reg, cmsb_reg, so_reg,
    f0_bus_stat_reg, f0_blk_stat_reg, f1_bus_stat_reg, f1_blk_stat_reg);
    input		reset;
    input		clk;
    input	[02:00]	cs_addr;
    input		route_si;
    input		route_ci;
    input		f0_load;
    input		f1_load;
    input		d0_load;
    input		d1_load;
    output	[01:00]	ce0;
    output	[01:00]	cl0;
    output	[01:00]	z0;
    output	[01:00]	ff0;
    output	[01:00]	ce1;
    output	[01:00]	cl1;
    output	[01:00]	z1;
    output	[01:00]	ff1;
    output	[01:00]	ov_msb;
    output	[01:00]	co_msb;
    output	[01:00]	cmsb;
    output	[01:00]	so;
    output	[01:00]	f0_bus_stat;
    output	[01:00]	f0_blk_stat;
    output	[01:00]	f1_bus_stat;
    output	[01:00]	f1_blk_stat;
    output	[01:00]	ce0_reg;
    output	[01:00]	cl0_reg;
    output	[01:00]	z0_reg;
    output	[01:00]	ff0_reg;
    output	[01:00]	ce1_reg;
    output	[01:00]	cl1_reg;
    output	[01:00]	z1_reg;
    output	[01:00]	ff1_reg;
    output	[01:00]	ov_msb_reg;
    output	[01:00]	co_msb_reg;
    output	[01:00]	cmsb_reg;
    output	[01:00]	so_reg;
    output	[01:00]	f0_bus_stat_reg;
    output	[01:00]	f0_blk_stat_reg;
    output	[01:00]	f1_bus_stat_reg;
    output	[01:00]	f1_blk_stat_reg;

    parameter	[207:0] cy_dpconfig_a	= {128'h0,32'hFF00_FFFF,48'h0};
    parameter	[07:00] d0_init_a	= 8'b0;
    parameter	[07:00] d1_init_a	= 8'b0;
    parameter	[07:00] a0_init_a	= 8'b0;
    parameter	[07:00] a1_init_a	= 8'b0;
    parameter	[207:0] cy_dpconfig_b	= {128'h0,32'hFF00_FFFF,48'h0};
    parameter	[07:00] d0_init_b	= 8'b0;
    parameter	[07:00] d1_init_b	= 8'b0;
    parameter	[07:00] a0_init_b	= 8'b0;
    parameter	[07:00] a1_init_b	= 8'b0;
    parameter	[01:00]	ce0_sync	= 2'b11;
    parameter	[01:00]	cl0_sync	= 2'b11;
    parameter	[01:00]	z0_sync		= 2'b11;
    parameter	[01:00]	ff0_sync	= 2'b11;
    parameter	[01:00]	ce1_sync	= 2'b11;
    parameter	[01:00]	cl1_sync	= 2'b11;
    parameter	[01:00]	z1_sync		= 2'b11;
    parameter	[01:00]	ff1_sync	= 2'b11;
    parameter	[01:00]	ov_msb_sync	= 2'b11;
    parameter	[01:00]	co_msb_sync	= 2'b11;
    parameter	[01:00]	cmsb_sync	= 2'b11;
    parameter	[01:00]	so_sync		= 2'b11;
    parameter	[01:00]	f0_bus_sync	= 2'b11;
    parameter	[01:00]	f0_blk_sync	= 2'b11;
    parameter	[01:00]	f1_bus_sync	= 2'b11;
    parameter	[01:00]	f1_blk_sync	= 2'b11;

    wire		carry, sh_right, sh_left, msb, cfb;
    wire	[01:00]	cmp_eq, cmp_lt, cmp_zero, cmp_ff, cap;

    defparam U0.cy_dpconfig	= cy_dpconfig_a;
    defparam U0.d0_init		= d0_init_a;
    defparam U0.d1_init		= d1_init_a;
    defparam U0.a0_init		= a0_init_a;
    defparam U0.a1_init		= a1_init_a;
    defparam U0.ce0_sync	= ce0_sync[0];
    defparam U0.cl0_sync	= cl0_sync[0];
    defparam U0.z0_sync		= z0_sync[0];
    defparam U0.ff0_sync	= ff0_sync[0];
    defparam U0.ce1_sync	= ce1_sync[0];
    defparam U0.cl1_sync	= cl1_sync[0];
    defparam U0.z1_sync		= z1_sync[0];
    defparam U0.ff1_sync	= ff1_sync[0];
    defparam U0.ov_msb_sync	= ov_msb_sync[0];
    defparam U0.co_msb_sync	= co_msb_sync[0];
    defparam U0.cmsb_sync	= cmsb_sync[0];
    defparam U0.so_sync		= so_sync[0];
    defparam U0.f0_bus_sync	= f0_bus_sync[0];
    defparam U0.f0_blk_sync	= f0_blk_sync[0];
    defparam U0.f1_bus_sync	= f1_bus_sync[0];
    defparam U0.f1_blk_sync	= f1_blk_sync[0];
    cy_psoc3_dp U0 (
	.reset			(reset),
	.clk			(clk),
	.cs_addr		(cs_addr),
	.route_si		(route_si),
	.route_ci		(route_ci),
	.f0_load		(f0_load),
	.f1_load		(f1_load),
	.d0_load		(d0_load),
	.d1_load		(d1_load),
	.ce0			(ce0[00]),
	.cl0			(cl0[00]),
	.z0			(z0[00]),
	.ff0			(ff0[00]),
	.ce1			(ce1[00]),
	.cl1			(cl1[00]),
	.z1			(z1[00]),
	.ff1			(ff1[00]),
	.ov_msb			(ov_msb[00]),
	.co_msb			(co_msb[00]),
	.cmsb			(cmsb[00]),
	.so			(so[00]),
	.f0_bus_stat		(f0_bus_stat[00]),
	.f0_blk_stat		(f0_blk_stat[00]),
	.f1_bus_stat		(f1_bus_stat[00]),
	.f1_blk_stat		(f1_blk_stat[00]),
	.ce0_reg		(ce0_reg[00]),
	.cl0_reg		(cl0_reg[00]),
	.z0_reg			(z0_reg[00]),
	.ff0_reg		(ff0_reg[00]),
	.ce1_reg		(ce1_reg[00]),
	.cl1_reg		(cl1_reg[00]),
	.z1_reg			(z1_reg[00]),
	.ff1_reg		(ff1_reg[00]),
	.ov_msb_reg		(ov_msb_reg[00]),
	.co_msb_reg		(co_msb_reg[00]),
	.cmsb_reg		(cmsb_reg[00]),
	.so_reg			(so_reg[00]),
	.f0_bus_stat_reg	(f0_bus_stat_reg[00]),
	.f0_blk_stat_reg	(f0_blk_stat_reg[00]),
	.f1_bus_stat_reg	(f1_bus_stat_reg[00]),
	.f1_blk_stat_reg	(f1_blk_stat_reg[00]),
	.ci			(1'b0),
	.co			(carry),
	.sir			(1'b0),
	.sor			(),
	.sil			(sh_right),
	.sol			(sh_left),
	.msbi			(msb),
	.msbo			(),
	.cei			(2'b00),
	.ceo			(cmp_eq),
	.cli			(2'b00),
	.clo			(cmp_lt),
	.zi			(2'b00),
	.zo			(cmp_zero),
	.fi			(2'b00),
	.fo			(cmp_ff),
	.capi			(2'b00),
	.capo			(cap),
	.cfbi			(1'b1),
	.cfbo			(cfb),
	.pi			(8'b00000000),
	.po			());

    defparam U1.cy_dpconfig	= cy_dpconfig_b;
    defparam U1.d0_init		= d0_init_b;
    defparam U1.d1_init		= d1_init_b;
    defparam U1.a0_init		= a0_init_b;
    defparam U1.a1_init		= a1_init_b;
    defparam U1.ce0_sync	= ce0_sync[1];
    defparam U1.cl0_sync	= cl0_sync[1];
    defparam U1.z0_sync		= z0_sync[1];
    defparam U1.ff0_sync	= ff0_sync[1];
    defparam U1.ce1_sync	= ce1_sync[1];
    defparam U1.cl1_sync	= cl1_sync[1];
    defparam U1.z1_sync		= z1_sync[1];
    defparam U1.ff1_sync	= ff1_sync[1];
    defparam U1.ov_msb_sync	= ov_msb_sync[1];
    defparam U1.co_msb_sync	= co_msb_sync[1];
    defparam U1.cmsb_sync	= cmsb_sync[1];
    defparam U1.so_sync		= so_sync[1];
    defparam U1.f0_bus_sync	= f0_bus_sync[1];
    defparam U1.f0_blk_sync	= f0_blk_sync[1];
    defparam U1.f1_bus_sync	= f1_bus_sync[1];
    defparam U1.f1_blk_sync	= f1_blk_sync[1];
    cy_psoc3_dp U1 		(
	.reset			(reset),
	.clk			(clk),
	.cs_addr		(cs_addr),
	.route_si		(route_si),
	.route_ci		(route_ci),
	.f0_load		(f0_load),
	.f1_load		(f1_load),
	.d0_load		(d0_load),
	.d1_load		(d1_load),
	.ce0			(ce0[01]),
	.cl0			(cl0[01]),
	.z0			(z0[01]),
	.ff0			(ff0[01]),
	.ce1			(ce1[01]),
	.cl1			(cl1[01]),
	.z1			(z1[01]),
	.ff1			(ff1[01]),
	.ov_msb			(ov_msb[01]),
	.co_msb			(co_msb[01]),
	.cmsb			(cmsb[01]),
	.so			(so[01]),
	.f0_bus_stat		(f0_bus_stat[01]),
	.f0_blk_stat		(f0_blk_stat[01]),
	.f1_bus_stat		(f1_bus_stat[01]),
	.f1_blk_stat		(f1_blk_stat[01]),
	.ce0_reg		(ce0_reg[01]),
	.cl0_reg		(cl0_reg[01]),
	.z0_reg			(z0_reg[01]),
	.ff0_reg		(ff0_reg[01]),
	.ce1_reg		(ce1_reg[01]),
	.cl1_reg		(cl1_reg[01]),
	.z1_reg			(z1_reg[01]),
	.ff1_reg		(ff1_reg[01]),
	.ov_msb_reg		(ov_msb_reg[01]),
	.co_msb_reg		(co_msb_reg[01]),
	.cmsb_reg		(cmsb_reg[01]),
	.so_reg			(so_reg[01]),
	.f0_bus_stat_reg	(f0_bus_stat_reg[01]),
	.f0_blk_stat_reg	(f0_blk_stat_reg[01]),
	.f1_bus_stat_reg	(f1_bus_stat_reg[01]),
	.f1_blk_stat_reg	(f1_blk_stat_reg[01]),
	.ci			(carry),
	.co			(),
	.sir			(sh_left),
	.sor			(sh_right),
	.sil			(1'b0),
	.sol			(),
	.msbi			(1'b0),
	.msbo			(msb),
	.cei			(cmp_eq),
	.ceo			(),
	.cli			(cmp_lt),
	.clo			(),
	.zi			(cmp_zero),
	.zo			(),
	.fi			(cmp_ff),
	.fo			(),
	.capi			(cap),
	.capo			(),
	.cfbi			(cfb),
	.cfbo			(),
	.pi			(8'b00000000),
	.po			());
endmodule

//
//	cy_psoc3_dp24
//

module cy_psoc3_dp24 (reset, clk,
    cs_addr, route_si, route_ci, f0_load, f1_load, d0_load, d1_load,
    ce0, cl0, z0, ff0, ce1, cl1, z1, ff1, ov_msb, co_msb, cmsb, so,
    f0_bus_stat, f0_blk_stat, f1_bus_stat, f1_blk_stat,
    ce0_reg, cl0_reg, z0_reg, ff0_reg, ce1_reg, cl1_reg, z1_reg,
    ff1_reg, ov_msb_reg, co_msb_reg, cmsb_reg, so_reg,
    f0_bus_stat_reg, f0_blk_stat_reg, f1_bus_stat_reg, f1_blk_stat_reg);
    input		reset;
    input		clk;
    input	[02:00]	cs_addr;
    input		route_si;
    input		route_ci;
    input		f0_load;
    input		f1_load;
    input		d0_load;
    input		d1_load;
    output	[02:00]	ce0;
    output	[02:00]	cl0;
    output	[02:00]	z0;
    output	[02:00]	ff0;
    output	[02:00]	ce1;
    output	[02:00]	cl1;
    output	[02:00]	z1;
    output	[02:00]	ff1;
    output	[02:00]	ov_msb;
    output	[02:00]	co_msb;
    output	[02:00]	cmsb;
    output	[02:00]	so;
    output	[02:00]	f0_bus_stat;
    output	[02:00]	f0_blk_stat;
    output	[02:00]	f1_bus_stat;
    output	[02:00]	f1_blk_stat;
    output	[02:00]	ce0_reg;
    output	[02:00]	cl0_reg;
    output	[02:00]	z0_reg;
    output	[02:00]	ff0_reg;
    output	[02:00]	ce1_reg;
    output	[02:00]	cl1_reg;
    output	[02:00]	z1_reg;
    output	[02:00]	ff1_reg;
    output	[02:00]	ov_msb_reg;
    output	[02:00]	co_msb_reg;
    output	[02:00]	cmsb_reg;
    output	[02:00]	so_reg;
    output	[02:00]	f0_bus_stat_reg;
    output	[02:00]	f0_blk_stat_reg;
    output	[02:00]	f1_bus_stat_reg;
    output	[02:00]	f1_blk_stat_reg;

    parameter	[207:0] cy_dpconfig_a	= {128'h0,32'hFF00_FFFF,48'h0};
    parameter	[07:00] d0_init_a	= 8'b0;
    parameter	[07:00] d1_init_a	= 8'b0;
    parameter	[07:00] a0_init_a	= 8'b0;
    parameter	[07:00] a1_init_a	= 8'b0;
    parameter	[207:0] cy_dpconfig_b	= {128'h0,32'hFF00_FFFF,48'h0};
    parameter	[07:00] d0_init_b	= 8'b0;
    parameter	[07:00] d1_init_b	= 8'b0;
    parameter	[07:00] a0_init_b	= 8'b0;
    parameter	[07:00] a1_init_b	= 8'b0;
    parameter	[207:0] cy_dpconfig_c	= {128'h0,32'hFF00_FFFF,48'h0};
    parameter	[07:00] d0_init_c	= 8'b0;
    parameter	[07:00] d1_init_c	= 8'b0;
    parameter	[07:00] a0_init_c	= 8'b0;
    parameter	[07:00] a1_init_c	= 8'b0;
    parameter	[02:00]	ce0_sync	= 3'b111;
    parameter	[02:00]	cl0_sync	= 3'b111;
    parameter	[02:00]	z0_sync		= 3'b111;
    parameter	[02:00]	ff0_sync	= 3'b111;
    parameter	[02:00]	ce1_sync	= 3'b111;
    parameter	[02:00]	cl1_sync	= 3'b111;
    parameter	[02:00]	z1_sync		= 3'b111;
    parameter	[02:00]	ff1_sync	= 3'b111;
    parameter	[02:00]	ov_msb_sync	= 3'b111;
    parameter	[02:00]	co_msb_sync	= 3'b111;
    parameter	[02:00]	cmsb_sync	= 3'b111;
    parameter	[02:00]	so_sync		= 3'b111;
    parameter	[02:00]	f0_bus_sync	= 3'b111;
    parameter	[02:00]	f0_blk_sync	= 3'b111;
    parameter	[02:00]	f1_bus_sync	= 3'b111;
    parameter	[02:00]	f1_blk_sync	= 3'b111;

    wire		carry0, sh_right0, sh_left0, msb0, cfb0;
    wire		carry1, sh_right1, sh_left1, msb1, cfb1;
    wire	[01:00]	cmp_eq0, cmp_lt0, cmp_zero0, cmp_ff0, cap0;
    wire	[01:00]	cmp_eq1, cmp_lt1, cmp_zero1, cmp_ff1, cap1;

    defparam U0.cy_dpconfig	= cy_dpconfig_a;
    defparam U0.d0_init		= d0_init_a;
    defparam U0.d1_init		= d1_init_a;
    defparam U0.a0_init		= a0_init_a;
    defparam U0.a1_init		= a1_init_a;
    defparam U0.ce0_sync	= ce0_sync[0];
    defparam U0.cl0_sync	= cl0_sync[0];
    defparam U0.z0_sync		= z0_sync[0];
    defparam U0.ff0_sync	= ff0_sync[0];
    defparam U0.ce1_sync	= ce1_sync[0];
    defparam U0.cl1_sync	= cl1_sync[0];
    defparam U0.z1_sync		= z1_sync[0];
    defparam U0.ff1_sync	= ff1_sync[0];
    defparam U0.ov_msb_sync	= ov_msb_sync[0];
    defparam U0.co_msb_sync	= co_msb_sync[0];
    defparam U0.cmsb_sync	= cmsb_sync[0];
    defparam U0.so_sync		= so_sync[0];
    defparam U0.f0_bus_sync	= f0_bus_sync[0];
    defparam U0.f0_blk_sync	= f0_blk_sync[0];
    defparam U0.f1_bus_sync	= f1_bus_sync[0];
    defparam U0.f1_blk_sync	= f1_blk_sync[0];
    cy_psoc3_dp U0 (
	.reset			(reset),
	.clk			(clk),
	.cs_addr		(cs_addr),
	.route_si		(route_si),
	.route_ci		(route_ci),
	.f0_load		(f0_load),
	.f1_load		(f1_load),
	.d0_load		(d0_load),
	.d1_load		(d1_load),
	.ce0			(ce0[00]),
	.cl0			(cl0[00]),
	.z0			(z0[00]),
	.ff0			(ff0[00]),
	.ce1			(ce1[00]),
	.cl1			(cl1[00]),
	.z1			(z1[00]),
	.ff1			(ff1[00]),
	.ov_msb			(ov_msb[00]),
	.co_msb			(co_msb[00]),
	.cmsb			(cmsb[00]),
	.so			(so[00]),
	.f0_bus_stat		(f0_bus_stat[00]),
	.f0_blk_stat		(f0_blk_stat[00]),
	.f1_bus_stat		(f1_bus_stat[00]),
	.f1_blk_stat		(f1_blk_stat[00]),
	.ce0_reg		(ce0_reg[00]),
	.cl0_reg		(cl0_reg[00]),
	.z0_reg			(z0_reg[00]),
	.ff0_reg		(ff0_reg[00]),
	.ce1_reg		(ce1_reg[00]),
	.cl1_reg		(cl1_reg[00]),
	.z1_reg			(z1_reg[00]),
	.ff1_reg		(ff1_reg[00]),
	.ov_msb_reg		(ov_msb_reg[00]),
	.co_msb_reg		(co_msb_reg[00]),
	.cmsb_reg		(cmsb_reg[00]),
	.so_reg			(so_reg[00]),
	.f0_bus_stat_reg	(f0_bus_stat_reg[00]),
	.f0_blk_stat_reg	(f0_blk_stat_reg[00]),
	.f1_bus_stat_reg	(f1_bus_stat_reg[00]),
	.f1_blk_stat_reg	(f1_blk_stat_reg[00]),
	.ci			(1'b0),
	.co			(carry0),
	.sir			(1'b0),
	.sor			(),
	.sil			(sh_right0),
	.sol			(sh_left0),
	.msbi			(msb0),
	.msbo			(),
	.cei			(2'b00),
	.ceo			(cmp_eq0),
	.cli			(2'b00),
	.clo			(cmp_lt0),
	.zi			(2'b00),
	.zo			(cmp_zero0),
	.fi			(2'b00),
	.fo			(cmp_ff0),
	.capi			(2'b00),
	.capo			(cap0),
	.cfbi			(1'b1),
	.cfbo			(cfb0),
	.pi			(8'b00000000),
	.po			());

    defparam U1.cy_dpconfig	= cy_dpconfig_b;
    defparam U1.d0_init		= d0_init_b;
    defparam U1.d1_init		= d1_init_b;
    defparam U1.a0_init		= a0_init_b;
    defparam U1.a1_init		= a1_init_b;
    defparam U1.ce0_sync	= ce0_sync[1];
    defparam U1.cl0_sync	= cl0_sync[1];
    defparam U1.z0_sync		= z0_sync[1];
    defparam U1.ff0_sync	= ff0_sync[1];
    defparam U1.ce1_sync	= ce1_sync[1];
    defparam U1.cl1_sync	= cl1_sync[1];
    defparam U1.z1_sync		= z1_sync[1];
    defparam U1.ff1_sync	= ff1_sync[1];
    defparam U1.ov_msb_sync	= ov_msb_sync[1];
    defparam U1.co_msb_sync	= co_msb_sync[1];
    defparam U1.cmsb_sync	= cmsb_sync[1];
    defparam U1.so_sync		= so_sync[1];
    defparam U1.f0_bus_sync	= f0_bus_sync[1];
    defparam U1.f0_blk_sync	= f0_blk_sync[1];
    defparam U1.f1_bus_sync	= f1_bus_sync[1];
    defparam U1.f1_blk_sync	= f1_blk_sync[1];
    cy_psoc3_dp U1 (
	.reset			(reset),
	.clk			(clk),
	.cs_addr		(cs_addr),
	.route_si		(route_si),
	.route_ci		(route_ci),
	.f0_load		(f0_load),
	.f1_load		(f1_load),
	.d0_load		(d0_load),
	.d1_load		(d1_load),
	.ce0			(ce0[01]),
	.cl0			(cl0[01]),
	.z0			(z0[01]),
	.ff0			(ff0[01]),
	.ce1			(ce1[01]),
	.cl1			(cl1[01]),
	.z1			(z1[01]),
	.ff1			(ff1[01]),
	.ov_msb			(ov_msb[01]),
	.co_msb			(co_msb[01]),
	.cmsb			(cmsb[01]),
	.so			(so[01]),
	.f0_bus_stat		(f0_bus_stat[01]),
	.f0_blk_stat		(f0_blk_stat[01]),
	.f1_bus_stat		(f1_bus_stat[01]),
	.f1_blk_stat		(f1_blk_stat[01]),
	.ce0_reg		(ce0_reg[01]),
	.cl0_reg		(cl0_reg[01]),
	.z0_reg			(z0_reg[01]),
	.ff0_reg		(ff0_reg[01]),
	.ce1_reg		(ce1_reg[01]),
	.cl1_reg		(cl1_reg[01]),
	.z1_reg			(z1_reg[01]),
	.ff1_reg		(ff1_reg[01]),
	.ov_msb_reg		(ov_msb_reg[01]),
	.co_msb_reg		(co_msb_reg[01]),
	.cmsb_reg		(cmsb_reg[01]),
	.so_reg			(so_reg[01]),
	.f0_bus_stat_reg	(f0_bus_stat_reg[01]),
	.f0_blk_stat_reg	(f0_blk_stat_reg[01]),
	.f1_bus_stat_reg	(f1_bus_stat_reg[01]),
	.f1_blk_stat_reg	(f1_blk_stat_reg[01]),
	.ci			(carry0),
	.co			(carry1),
	.sir			(sh_left0),
	.sor			(sh_right0),
	.sil			(sh_right1),
	.sol			(sh_left1),
	.msbi			(msb1),
	.msbo			(msb0),
	.cei			(cmp_eq0),
	.ceo			(cmp_eq1),
	.cli			(cmp_lt0),
	.clo			(cmp_lt1),
	.zi			(cmp_zero0),
	.zo			(cmp_zero1),
	.fi			(cmp_ff0),
	.fo			(cmp_ff1),
	.capi			(cap0),
	.capo			(cap1),
	.cfbi			(cfb0),
	.cfbo			(cfb1),
	.pi			(8'b00000000),
	.po			());

    defparam U2.cy_dpconfig	= cy_dpconfig_c;
    defparam U2.d0_init		= d0_init_c;
    defparam U2.d1_init		= d1_init_c;
    defparam U2.a0_init		= a0_init_c;
    defparam U2.a1_init		= a1_init_c;
    defparam U2.ce0_sync	= ce0_sync[2];
    defparam U2.cl0_sync	= cl0_sync[2];
    defparam U2.z0_sync		= z0_sync[2];
    defparam U2.ff0_sync	= ff0_sync[2];
    defparam U2.ce1_sync	= ce1_sync[2];
    defparam U2.cl1_sync	= cl1_sync[2];
    defparam U2.z1_sync		= z1_sync[2];
    defparam U2.ff1_sync	= ff1_sync[2];
    defparam U2.ov_msb_sync	= ov_msb_sync[2];
    defparam U2.co_msb_sync	= co_msb_sync[2];
    defparam U2.cmsb_sync	= cmsb_sync[2];
    defparam U2.so_sync		= so_sync[2];
    defparam U2.f0_bus_sync	= f0_bus_sync[2];
    defparam U2.f0_blk_sync	= f0_blk_sync[2];
    defparam U2.f1_bus_sync	= f1_bus_sync[2];
    defparam U2.f1_blk_sync	= f1_blk_sync[2];
    cy_psoc3_dp U2 (
	.reset			(reset),
	.clk			(clk),
	.cs_addr		(cs_addr),
	.route_si		(route_si),
	.route_ci		(route_ci),
	.f0_load		(f0_load),
	.f1_load		(f1_load),
	.d0_load		(d0_load),
	.d1_load		(d1_load),
	.ce0			(ce0[02]),
	.cl0			(cl0[02]),
	.z0			(z0[02]),
	.ff0			(ff0[02]),
	.ce1			(ce1[02]),
	.cl1			(cl1[02]),
	.z1			(z1[02]),
	.ff1			(ff1[02]),
	.ov_msb			(ov_msb[02]),
	.co_msb			(co_msb[02]),
	.cmsb			(cmsb[02]),
	.so			(so[02]),
	.f0_bus_stat		(f0_bus_stat[02]),
	.f0_blk_stat		(f0_blk_stat[02]),
	.f1_bus_stat		(f1_bus_stat[02]),
	.f1_blk_stat		(f1_blk_stat[02]),
	.ce0_reg		(ce0_reg[02]),
	.cl0_reg		(cl0_reg[02]),
	.z0_reg			(z0_reg[02]),
	.ff0_reg		(ff0_reg[02]),
	.ce1_reg		(ce1_reg[02]),
	.cl1_reg		(cl1_reg[02]),
	.z1_reg			(z1_reg[02]),
	.ff1_reg		(ff1_reg[02]),
	.ov_msb_reg		(ov_msb_reg[02]),
	.co_msb_reg		(co_msb_reg[02]),
	.cmsb_reg		(cmsb_reg[02]),
	.so_reg			(so_reg[02]),
	.f0_bus_stat_reg	(f0_bus_stat_reg[02]),
	.f0_blk_stat_reg	(f0_blk_stat_reg[02]),
	.f1_bus_stat_reg	(f1_bus_stat_reg[02]),
	.f1_blk_stat_reg	(f1_blk_stat_reg[02]),
	.ci			(carry1),
	.co			(),
	.sir			(sh_left1),
	.sor			(sh_right1),
	.sil			(1'b0),
	.sol			(),
	.msbi			(1'b0),
	.msbo			(msb1),
	.cei			(cmp_eq1),
	.ceo			(),
	.cli			(cmp_lt1),
	.clo			(),
	.zi			(cmp_zero1),
	.zo			(),
	.fi			(cmp_ff1),
	.fo			(),
	.capi			(cap1),
	.capo			(),
	.cfbi			(cfb1),
	.cfbo			(),
	.pi			(8'b00000000),
	.po			());
endmodule

//
//	cy_psoc3_dp32
//

module cy_psoc3_dp32 (reset, clk,
    cs_addr, route_si, route_ci, f0_load, f1_load, d0_load, d1_load,
    ce0, cl0, z0, ff0, ce1, cl1, z1, ff1, ov_msb, co_msb, cmsb, so,
    f0_bus_stat, f0_blk_stat, f1_bus_stat, f1_blk_stat,
    ce0_reg, cl0_reg, z0_reg, ff0_reg, ce1_reg, cl1_reg, z1_reg,
    ff1_reg, ov_msb_reg, co_msb_reg, cmsb_reg, so_reg,
    f0_bus_stat_reg, f0_blk_stat_reg, f1_bus_stat_reg, f1_blk_stat_reg);
    input		reset;
    input		clk;
    input	[02:00]	cs_addr;
    input		route_si;
    input		route_ci;
    input		f0_load;
    input		f1_load;
    input		d0_load;
    input		d1_load;
    output	[03:00]	ce0;
    output	[03:00]	cl0;
    output	[03:00]	z0;
    output	[03:00]	ff0;
    output	[03:00]	ce1;
    output	[03:00]	cl1;
    output	[03:00]	z1;
    output	[03:00]	ff1;
    output	[03:00]	ov_msb;
    output	[03:00]	co_msb;
    output	[03:00]	cmsb;
    output	[03:00]	so;
    output	[03:00]	f0_bus_stat;
    output	[03:00]	f0_blk_stat;
    output	[03:00]	f1_bus_stat;
    output	[03:00]	f1_blk_stat;
    output	[03:00]	ce0_reg;
    output	[03:00]	cl0_reg;
    output	[03:00]	z0_reg;
    output	[03:00]	ff0_reg;
    output	[03:00]	ce1_reg;
    output	[03:00]	cl1_reg;
    output	[03:00]	z1_reg;
    output	[03:00]	ff1_reg;
    output	[03:00]	ov_msb_reg;
    output	[03:00]	co_msb_reg;
    output	[03:00]	cmsb_reg;
    output	[03:00]	so_reg;
    output	[03:00]	f0_bus_stat_reg;
    output	[03:00]	f0_blk_stat_reg;
    output	[03:00]	f1_bus_stat_reg;
    output	[03:00]	f1_blk_stat_reg;

    parameter	[207:0] cy_dpconfig_a	= {128'h0,32'hFF00_FFFF,48'h0};
    parameter	[07:00] d0_init_a	= 8'b0;
    parameter	[07:00] d1_init_a	= 8'b0;
    parameter	[07:00] a0_init_a	= 8'b0;
    parameter	[07:00] a1_init_a	= 8'b0;
    parameter	[207:0] cy_dpconfig_b	= {128'h0,32'hFF00_FFFF,48'h0};
    parameter	[07:00] d0_init_b	= 8'b0;
    parameter	[07:00] d1_init_b	= 8'b0;
    parameter	[07:00] a0_init_b	= 8'b0;
    parameter	[07:00] a1_init_b	= 8'b0;
    parameter	[207:0] cy_dpconfig_c	= {128'h0,32'hFF00_FFFF,48'h0};
    parameter	[07:00] d0_init_c	= 8'b0;
    parameter	[07:00] d1_init_c	= 8'b0;
    parameter	[07:00] a0_init_c	= 8'b0;
    parameter	[07:00] a1_init_c	= 8'b0;
    parameter	[207:0] cy_dpconfig_d	= {128'h0,32'hFF00_FFFF,48'h0};
    parameter	[07:00] d0_init_d	= 8'b0;
    parameter	[07:00] d1_init_d	= 8'b0;
    parameter	[07:00] a0_init_d	= 8'b0;
    parameter	[07:00] a1_init_d	= 8'b0;
    parameter	[03:00]	ce0_sync	= 4'b1111;
    parameter	[03:00]	cl0_sync	= 4'b1111;
    parameter	[03:00]	z0_sync		= 4'b1111;
    parameter	[03:00]	ff0_sync	= 4'b1111;
    parameter	[03:00]	ce1_sync	= 4'b1111;
    parameter	[03:00]	cl1_sync	= 4'b1111;
    parameter	[03:00]	z1_sync		= 4'b1111;
    parameter	[03:00]	ff1_sync	= 4'b1111;
    parameter	[03:00]	ov_msb_sync	= 4'b1111;
    parameter	[03:00]	co_msb_sync	= 4'b1111;
    parameter	[03:00]	cmsb_sync	= 4'b1111;
    parameter	[03:00]	so_sync		= 4'b1111;
    parameter	[03:00]	f0_bus_sync	= 4'b1111;
    parameter	[03:00]	f0_blk_sync	= 4'b1111;
    parameter	[03:00]	f1_bus_sync	= 4'b1111;
    parameter	[03:00]	f1_blk_sync	= 4'b1111;

    wire		carry0, sh_right0, sh_left0, msb0, cfb0;
    wire		carry1, sh_right1, sh_left1, msb1, cfb1;
    wire		carry2, sh_right2, sh_left2, msb2, cfb2;
    wire	[01:00]	cmp_eq0, cmp_lt0, cmp_zero0, cmp_ff0, cap0;
    wire	[01:00]	cmp_eq1, cmp_lt1, cmp_zero1, cmp_ff1, cap1;
    wire	[01:00]	cmp_eq2, cmp_lt2, cmp_zero2, cmp_ff2, cap2;

    defparam U0.cy_dpconfig	= cy_dpconfig_a;
    defparam U0.d0_init		= d0_init_a;
    defparam U0.d1_init		= d1_init_a;
    defparam U0.a0_init		= a0_init_a;
    defparam U0.a1_init		= a1_init_a;
    defparam U0.ce0_sync	= ce0_sync[0];
    defparam U0.cl0_sync	= cl0_sync[0];
    defparam U0.z0_sync		= z0_sync[0];
    defparam U0.ff0_sync	= ff0_sync[0];
    defparam U0.ce1_sync	= ce1_sync[0];
    defparam U0.cl1_sync	= cl1_sync[0];
    defparam U0.z1_sync		= z1_sync[0];
    defparam U0.ff1_sync	= ff1_sync[0];
    defparam U0.ov_msb_sync	= ov_msb_sync[0];
    defparam U0.co_msb_sync	= co_msb_sync[0];
    defparam U0.cmsb_sync	= cmsb_sync[0];
    defparam U0.so_sync		= so_sync[0];
    defparam U0.f0_bus_sync	= f0_bus_sync[0];
    defparam U0.f0_blk_sync	= f0_blk_sync[0];
    defparam U0.f1_bus_sync	= f1_bus_sync[0];
    defparam U0.f1_blk_sync	= f1_blk_sync[0];
    cy_psoc3_dp U0 (
	.reset			(reset),
	.clk			(clk),
	.cs_addr		(cs_addr),
	.route_si		(route_si),
	.route_ci		(route_ci),
	.f0_load		(f0_load),
	.f1_load		(f1_load),
	.d0_load		(d0_load),
	.d1_load		(d1_load),
	.ce0			(ce0[00]),
	.cl0			(cl0[00]),
	.z0			(z0[00]),
	.ff0			(ff0[00]),
	.ce1			(ce1[00]),
	.cl1			(cl1[00]),
	.z1			(z1[00]),
	.ff1			(ff1[00]),
	.ov_msb			(ov_msb[00]),
	.co_msb			(co_msb[00]),
	.cmsb			(cmsb[00]),
	.so			(so[00]),
	.f0_bus_stat		(f0_bus_stat[00]),
	.f0_blk_stat		(f0_blk_stat[00]),
	.f1_bus_stat		(f1_bus_stat[00]),
	.f1_blk_stat		(f1_blk_stat[00]),
	.ce0_reg		(ce0_reg[00]),
	.cl0_reg		(cl0_reg[00]),
	.z0_reg			(z0_reg[00]),
	.ff0_reg		(ff0_reg[00]),
	.ce1_reg		(ce1_reg[00]),
	.cl1_reg		(cl1_reg[00]),
	.z1_reg			(z1_reg[00]),
	.ff1_reg		(ff1_reg[00]),
	.ov_msb_reg		(ov_msb_reg[00]),
	.co_msb_reg		(co_msb_reg[00]),
	.cmsb_reg		(cmsb_reg[00]),
	.so_reg			(so_reg[00]),
	.f0_bus_stat_reg	(f0_bus_stat_reg[00]),
	.f0_blk_stat_reg	(f0_blk_stat_reg[00]),
	.f1_bus_stat_reg	(f1_bus_stat_reg[00]),
	.f1_blk_stat_reg	(f1_blk_stat_reg[00]),
	.ci			(1'b0),
	.co			(carry0),
	.sir			(1'b0),
	.sor			(),
	.sil			(sh_right0),
	.sol			(sh_left0),
	.msbi			(msb0),
	.msbo			(),
	.cei			(2'b00),
	.ceo			(cmp_eq0),
	.cli			(2'b00),
	.clo			(cmp_lt0),
	.zi			(2'b00),
	.zo			(cmp_zero0),
	.fi			(2'b00),
	.fo			(cmp_ff0),
	.capi			(2'b00),
	.capo			(cap0),
	.cfbi			(1'b1),
	.cfbo			(cfb0),
	.pi			(8'b00000000),
	.po			());

    defparam U1.cy_dpconfig	= cy_dpconfig_b;
    defparam U1.d0_init		= d0_init_b;
    defparam U1.d1_init		= d1_init_b;
    defparam U1.a0_init		= a0_init_b;
    defparam U1.a1_init		= a1_init_b;
    defparam U1.ce0_sync	= ce0_sync[1];
    defparam U1.cl0_sync	= cl0_sync[1];
    defparam U1.z0_sync		= z0_sync[1];
    defparam U1.ff0_sync	= ff0_sync[1];
    defparam U1.ce1_sync	= ce1_sync[1];
    defparam U1.cl1_sync	= cl1_sync[1];
    defparam U1.z1_sync		= z1_sync[1];
    defparam U1.ff1_sync	= ff1_sync[1];
    defparam U1.ov_msb_sync	= ov_msb_sync[1];
    defparam U1.co_msb_sync	= co_msb_sync[1];
    defparam U1.cmsb_sync	= cmsb_sync[1];
    defparam U1.so_sync		= so_sync[1];
    defparam U1.f0_bus_sync	= f0_bus_sync[1];
    defparam U1.f0_blk_sync	= f0_blk_sync[1];
    defparam U1.f1_bus_sync	= f1_bus_sync[1];
    defparam U1.f1_blk_sync	= f1_blk_sync[1];
    cy_psoc3_dp U1 (
	.reset			(reset),
	.clk			(clk),
	.cs_addr		(cs_addr),
	.route_si		(route_si),
	.route_ci		(route_ci),
	.f0_load		(f0_load),
	.f1_load		(f1_load),
	.d0_load		(d0_load),
	.d1_load		(d1_load),
	.ce0			(ce0[01]),
	.cl0			(cl0[01]),
	.z0			(z0[01]),
	.ff0			(ff0[01]),
	.ce1			(ce1[01]),
	.cl1			(cl1[01]),
	.z1			(z1[01]),
	.ff1			(ff1[01]),
	.ov_msb			(ov_msb[01]),
	.co_msb			(co_msb[01]),
	.cmsb			(cmsb[01]),
	.so			(so[01]),
	.f0_bus_stat		(f0_bus_stat[01]),
	.f0_blk_stat		(f0_blk_stat[01]),
	.f1_bus_stat		(f1_bus_stat[01]),
	.f1_blk_stat		(f1_blk_stat[01]),
	.ce0_reg		(ce0_reg[01]),
	.cl0_reg		(cl0_reg[01]),
	.z0_reg			(z0_reg[01]),
	.ff0_reg		(ff0_reg[01]),
	.ce1_reg		(ce1_reg[01]),
	.cl1_reg		(cl1_reg[01]),
	.z1_reg			(z1_reg[01]),
	.ff1_reg		(ff1_reg[01]),
	.ov_msb_reg		(ov_msb_reg[01]),
	.co_msb_reg		(co_msb_reg[01]),
	.cmsb_reg		(cmsb_reg[01]),
	.so_reg			(so_reg[01]),
	.f0_bus_stat_reg	(f0_bus_stat_reg[01]),
	.f0_blk_stat_reg	(f0_blk_stat_reg[01]),
	.f1_bus_stat_reg	(f1_bus_stat_reg[01]),
	.f1_blk_stat_reg	(f1_blk_stat_reg[01]),
	.ci			(carry0),
	.co			(carry1),
	.sir			(sh_left0),
	.sor			(sh_right0),
	.sil			(sh_right1),
	.sol			(sh_left1),
	.msbi			(msb1),
	.msbo			(msb0),
	.cei			(cmp_eq0),
	.ceo			(cmp_eq1),
	.cli			(cmp_lt0),
	.clo			(cmp_lt1),
	.zi			(cmp_zero0),
	.zo			(cmp_zero1),
	.fi			(cmp_ff0),
	.fo			(cmp_ff1),
	.capi			(cap0),
	.capo			(cap1),
	.cfbi			(cfb0),
	.cfbo			(cfb1),
	.pi			(8'b00000000),
	.po			());

    defparam U2.cy_dpconfig	= cy_dpconfig_c;
    defparam U2.d0_init		= d0_init_c;
    defparam U2.d1_init		= d1_init_c;
    defparam U2.a0_init		= a0_init_c;
    defparam U2.a1_init		= a1_init_c;
    defparam U2.ce0_sync	= ce0_sync[2];
    defparam U2.cl0_sync	= cl0_sync[2];
    defparam U2.z0_sync		= z0_sync[2];
    defparam U2.ff0_sync	= ff0_sync[2];
    defparam U2.ce1_sync	= ce1_sync[2];
    defparam U2.cl1_sync	= cl1_sync[2];
    defparam U2.z1_sync		= z1_sync[2];
    defparam U2.ff1_sync	= ff1_sync[2];
    defparam U2.ov_msb_sync	= ov_msb_sync[2];
    defparam U2.co_msb_sync	= co_msb_sync[2];
    defparam U2.cmsb_sync	= cmsb_sync[2];
    defparam U2.so_sync		= so_sync[2];
    defparam U2.f0_bus_sync	= f0_bus_sync[2];
    defparam U2.f0_blk_sync	= f0_blk_sync[2];
    defparam U2.f1_bus_sync	= f1_bus_sync[2];
    defparam U2.f1_blk_sync	= f1_blk_sync[2];
    cy_psoc3_dp U2 (
	.reset			(reset),
	.clk			(clk),
	.cs_addr		(cs_addr),
	.route_si		(route_si),
	.route_ci		(route_ci),
	.f0_load		(f0_load),
	.f1_load		(f1_load),
	.d0_load		(d0_load),
	.d1_load		(d1_load),
	.ce0			(ce0[02]),
	.cl0			(cl0[02]),
	.z0			(z0[02]),
	.ff0			(ff0[02]),
	.ce1			(ce1[02]),
	.cl1			(cl1[02]),
	.z1			(z1[02]),
	.ff1			(ff1[02]),
	.ov_msb			(ov_msb[02]),
	.co_msb			(co_msb[02]),
	.cmsb			(cmsb[02]),
	.so			(so[02]),
	.f0_bus_stat		(f0_bus_stat[02]),
	.f0_blk_stat		(f0_blk_stat[02]),
	.f1_bus_stat		(f1_bus_stat[02]),
	.f1_blk_stat		(f1_blk_stat[02]),
	.ce0_reg		(ce0_reg[02]),
	.cl0_reg		(cl0_reg[02]),
	.z0_reg			(z0_reg[02]),
	.ff0_reg		(ff0_reg[02]),
	.ce1_reg		(ce1_reg[02]),
	.cl1_reg		(cl1_reg[02]),
	.z1_reg			(z1_reg[02]),
	.ff1_reg		(ff1_reg[02]),
	.ov_msb_reg		(ov_msb_reg[02]),
	.co_msb_reg		(co_msb_reg[02]),
	.cmsb_reg		(cmsb_reg[02]),
	.so_reg			(so_reg[02]),
	.f0_bus_stat_reg	(f0_bus_stat_reg[02]),
	.f0_blk_stat_reg	(f0_blk_stat_reg[02]),
	.f1_bus_stat_reg	(f1_bus_stat_reg[02]),
	.f1_blk_stat_reg	(f1_blk_stat_reg[02]),
	.ci			(carry1),
	.co			(carry2),
	.sir			(sh_left1),
	.sor			(sh_right1),
	.sil			(sh_right2),
	.sol			(sh_left2),
	.msbi			(msb2),
	.msbo			(msb1),
	.cei			(cmp_eq1),
	.ceo			(cmp_eq2),
	.cli			(cmp_lt1),
	.clo			(cmp_lt2),
	.zi			(cmp_zero1),
	.zo			(cmp_zero2),
	.fi			(cmp_ff1),
	.fo			(cmp_ff2),
	.capi			(cap1),
	.capo			(cap2),
	.cfbi			(cfb1),
	.cfbo			(cfb2),
	.pi			(8'b00000000),
	.po			());

    defparam U3.cy_dpconfig	= cy_dpconfig_d;
    defparam U3.d0_init		= d0_init_d;
    defparam U3.d1_init		= d1_init_d;
    defparam U3.a0_init		= a0_init_d;
    defparam U3.a1_init		= a1_init_d;
    defparam U3.ce0_sync	= ce0_sync[3];
    defparam U3.cl0_sync	= cl0_sync[3];
    defparam U3.z0_sync		= z0_sync[3];
    defparam U3.ff0_sync	= ff0_sync[3];
    defparam U3.ce1_sync	= ce1_sync[3];
    defparam U3.cl1_sync	= cl1_sync[3];
    defparam U3.z1_sync		= z1_sync[3];
    defparam U3.ff1_sync	= ff1_sync[3];
    defparam U3.ov_msb_sync	= ov_msb_sync[3];
    defparam U3.co_msb_sync	= co_msb_sync[3];
    defparam U3.cmsb_sync	= cmsb_sync[3];
    defparam U3.so_sync		= so_sync[3];
    defparam U3.f0_bus_sync	= f0_bus_sync[3];
    defparam U3.f0_blk_sync	= f0_blk_sync[3];
    defparam U3.f1_bus_sync	= f1_bus_sync[3];
    defparam U3.f1_blk_sync	= f1_blk_sync[3];
    cy_psoc3_dp U3 (
	.reset			(reset),
	.clk			(clk),
	.cs_addr		(cs_addr),
	.route_si		(route_si),
	.route_ci		(route_ci),
	.f0_load		(f0_load),
	.f1_load		(f1_load),
	.d0_load		(d0_load),
	.d1_load		(d1_load),
	.ce0			(ce0[03]),
	.cl0			(cl0[03]),
	.z0			(z0[03]),
	.ff0			(ff0[03]),
	.ce1			(ce1[03]),
	.cl1			(cl1[03]),
	.z1			(z1[03]),
	.ff1			(ff1[03]),
	.ov_msb			(ov_msb[03]),
	.co_msb			(co_msb[03]),
	.cmsb			(cmsb[03]),
	.so			(so[03]),
	.f0_bus_stat		(f0_bus_stat[03]),
	.f0_blk_stat		(f0_blk_stat[03]),
	.f1_bus_stat		(f1_bus_stat[03]),
	.f1_blk_stat		(f1_blk_stat[03]),
	.ce0_reg		(ce0_reg[03]),
	.cl0_reg		(cl0_reg[03]),
	.z0_reg			(z0_reg[03]),
	.ff0_reg		(ff0_reg[03]),
	.ce1_reg		(ce1_reg[03]),
	.cl1_reg		(cl1_reg[03]),
	.z1_reg			(z1_reg[03]),
	.ff1_reg		(ff1_reg[03]),
	.ov_msb_reg		(ov_msb_reg[03]),
	.co_msb_reg		(co_msb_reg[03]),
	.cmsb_reg		(cmsb_reg[03]),
	.so_reg			(so_reg[03]),
	.f0_bus_stat_reg	(f0_bus_stat_reg[03]),
	.f0_blk_stat_reg	(f0_blk_stat_reg[03]),
	.f1_bus_stat_reg	(f1_bus_stat_reg[03]),
	.f1_blk_stat_reg	(f1_blk_stat_reg[03]),
	.ci			(carry2),
	.co			(),
	.sir			(sh_left2),
	.sor			(sh_right2),
	.sil			(1'b0),
	.sol			(),
	.msbi			(1'b0),
	.msbo			(msb2),
	.cei			(cmp_eq2),
	.ceo			(),
	.cli			(cmp_lt2),
	.clo			(),
	.zi			(cmp_zero2),
	.zo			(),
	.fi			(cmp_ff2),
	.fo			(),
	.capi			(cap2),
	.capo			(),
	.cfbi			(cfb2),
	.cfbo			(),
	.pi			(8'b00000000),
	.po			());
endmodule

`endif
